-- Copyright 2002    Chuck Benz, Hollis, NH   
-- Copyright 2020    Frans Schreuder
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.


-- The information and description contained herein is the
-- property of Chuck Benz.
--
-- Permission is granted for any reuse of this information
-- and description as long as this copyright notice is
-- preserved.  Modifications may be made as long as this
-- notice is preserved.

-- Changelog:
-- 11 October  2002: Chuck Benz: updated with clearer messages, and checking decodeout
-- 3  November 2020: Frans Schreuder: Translated to VHDL, added UVVM testbench

library ieee;
use ieee.std_logic_1164.all;

package lookup_8b10b is

  type slv9_array is array(natural range <>) of std_logic_vector(8 downto 0);
  
  type code_type is record
    k : std_logic;
    val_8b : std_logic_vector(7 downto 0);
    val_10b_neg : std_logic_vector(9 downto 0);
    val_10b_pos : std_logic_vector(9 downto 0);
    disp_flip : std_logic;
  end record;
  
  type code_type_array is array(natural range <>) of code_type;
    

  constant code8b10b: code_type_array(0 to 267) := (
      ('0', "00000000", "1001110100", "0110001011", '0'),
      ('0', "00000001", "0111010100", "1000101011", '0'),
      ('0', "00000010", "1011010100", "0100101011", '0'),
      ('0', "00000011", "1100011011", "1100010100", '1'),
      ('0', "00000100", "1101010100", "0010101011", '0'),
      ('0', "00000101", "1010011011", "1010010100", '1'),
      ('0', "00000110", "0110011011", "0110010100", '1'),
      ('0', "00000111", "1110001011", "0001110100", '1'),
      ('0', "00001000", "1110010100", "0001101011", '0'),
      ('0', "00001001", "1001011011", "1001010100", '1'),
      ('0', "00001010", "0101011011", "0101010100", '1'),
      ('0', "00001011", "1101001011", "1101000100", '1'),
      ('0', "00001100", "0011011011", "0011010100", '1'),
      ('0', "00001101", "1011001011", "1011000100", '1'),
      ('0', "00001110", "0111001011", "0111000100", '1'),
      ('0', "00001111", "0101110100", "1010001011", '0'),
      ('0', "00010000", "0110110100", "1001001011", '0'),
      ('0', "00010001", "1000111011", "1000110100", '1'),
      ('0', "00010010", "0100111011", "0100110100", '1'),
      ('0', "00010011", "1100101011", "1100100100", '1'),
      ('0', "00010100", "0010111011", "0010110100", '1'),
      ('0', "00010101", "1010101011", "1010100100", '1'),
      ('0', "00010110", "0110101011", "0110100100", '1'),
      ('0', "00010111", "1110100100", "0001011011", '0'),
      ('0', "00011000", "1100110100", "0011001011", '0'),
      ('0', "00011001", "1001101011", "1001100100", '1'),
      ('0', "00011010", "0101101011", "0101100100", '1'),
      ('0', "00011011", "1101100100", "0010011011", '0'),
      ('0', "00011100", "0011101011", "0011100100", '1'),
      ('0', "00011101", "1011100100", "0100011011", '0'),
      ('0', "00011110", "0111100100", "1000011011", '0'),
      ('0', "00011111", "1010110100", "0101001011", '0'),
      ('0', "00100000", "1001111001", "0110001001", '1'),
      ('0', "00100001", "0111011001", "1000101001", '1'),
      ('0', "00100010", "1011011001", "0100101001", '1'),
      ('0', "00100011", "1100011001", "1100011001", '0'),
      ('0', "00100100", "1101011001", "0010101001", '1'),
      ('0', "00100101", "1010011001", "1010011001", '0'),
      ('0', "00100110", "0110011001", "0110011001", '0'),
      ('0', "00100111", "1110001001", "0001111001", '0'),
      ('0', "00101000", "1110011001", "0001101001", '1'),
      ('0', "00101001", "1001011001", "1001011001", '0'),
      ('0', "00101010", "0101011001", "0101011001", '0'),
      ('0', "00101011", "1101001001", "1101001001", '0'),
      ('0', "00101100", "0011011001", "0011011001", '0'),
      ('0', "00101101", "1011001001", "1011001001", '0'),
      ('0', "00101110", "0111001001", "0111001001", '0'),
      ('0', "00101111", "0101111001", "1010001001", '1'),
      ('0', "00110000", "0110111001", "1001001001", '1'),
      ('0', "00110001", "1000111001", "1000111001", '0'),
      ('0', "00110010", "0100111001", "0100111001", '0'),
      ('0', "00110011", "1100101001", "1100101001", '0'),
      ('0', "00110100", "0010111001", "0010111001", '0'),
      ('0', "00110101", "1010101001", "1010101001", '0'),
      ('0', "00110110", "0110101001", "0110101001", '0'),
      ('0', "00110111", "1110101001", "0001011001", '1'),
      ('0', "00111000", "1100111001", "0011001001", '1'),
      ('0', "00111001", "1001101001", "1001101001", '0'),
      ('0', "00111010", "0101101001", "0101101001", '0'),
      ('0', "00111011", "1101101001", "0010011001", '1'),
      ('0', "00111100", "0011101001", "0011101001", '0'),
      ('0', "00111101", "1011101001", "0100011001", '1'),
      ('0', "00111110", "0111101001", "1000011001", '1'),
      ('0', "00111111", "1010111001", "0101001001", '1'),
      ('0', "01000000", "1001110101", "0110000101", '1'),
      ('0', "01000001", "0111010101", "1000100101", '1'),
      ('0', "01000010", "1011010101", "0100100101", '1'),
      ('0', "01000011", "1100010101", "1100010101", '0'),
      ('0', "01000100", "1101010101", "0010100101", '1'),
      ('0', "01000101", "1010010101", "1010010101", '0'),
      ('0', "01000110", "0110010101", "0110010101", '0'),
      ('0', "01000111", "1110000101", "0001110101", '0'),
      ('0', "01001000", "1110010101", "0001100101", '1'),
      ('0', "01001001", "1001010101", "1001010101", '0'),
      ('0', "01001010", "0101010101", "0101010101", '0'),
      ('0', "01001011", "1101000101", "1101000101", '0'),
      ('0', "01001100", "0011010101", "0011010101", '0'),
      ('0', "01001101", "1011000101", "1011000101", '0'),
      ('0', "01001110", "0111000101", "0111000101", '0'),
      ('0', "01001111", "0101110101", "1010000101", '1'),
      ('0', "01010000", "0110110101", "1001000101", '1'),
      ('0', "01010001", "1000110101", "1000110101", '0'),
      ('0', "01010010", "0100110101", "0100110101", '0'),
      ('0', "01010011", "1100100101", "1100100101", '0'),
      ('0', "01010100", "0010110101", "0010110101", '0'),
      ('0', "01010101", "1010100101", "1010100101", '0'),
      ('0', "01010110", "0110100101", "0110100101", '0'),
      ('0', "01010111", "1110100101", "0001010101", '1'),
      ('0', "01011000", "1100110101", "0011000101", '1'),
      ('0', "01011001", "1001100101", "1001100101", '0'),
      ('0', "01011010", "0101100101", "0101100101", '0'),
      ('0', "01011011", "1101100101", "0010010101", '1'),
      ('0', "01011100", "0011100101", "0011100101", '0'),
      ('0', "01011101", "1011100101", "0100010101", '1'),
      ('0', "01011110", "0111100101", "1000010101", '1'),
      ('0', "01011111", "1010110101", "0101000101", '1'),
      ('0', "01100000", "1001110011", "0110001100", '1'),
      ('0', "01100001", "0111010011", "1000101100", '1'),
      ('0', "01100010", "1011010011", "0100101100", '1'),
      ('0', "01100011", "1100011100", "1100010011", '0'),
      ('0', "01100100", "1101010011", "0010101100", '1'),
      ('0', "01100101", "1010011100", "1010010011", '0'),
      ('0', "01100110", "0110011100", "0110010011", '0'),
      ('0', "01100111", "1110001100", "0001110011", '0'),
      ('0', "01101000", "1110010011", "0001101100", '1'),
      ('0', "01101001", "1001011100", "1001010011", '0'),
      ('0', "01101010", "0101011100", "0101010011", '0'),
      ('0', "01101011", "1101001100", "1101000011", '0'),
      ('0', "01101100", "0011011100", "0011010011", '0'),
      ('0', "01101101", "1011001100", "1011000011", '0'),
      ('0', "01101110", "0111001100", "0111000011", '0'),
      ('0', "01101111", "0101110011", "1010001100", '1'),
      ('0', "01110000", "0110110011", "1001001100", '1'),
      ('0', "01110001", "1000111100", "1000110011", '0'),
      ('0', "01110010", "0100111100", "0100110011", '0'),
      ('0', "01110011", "1100101100", "1100100011", '0'),
      ('0', "01110100", "0010111100", "0010110011", '0'),
      ('0', "01110101", "1010101100", "1010100011", '0'),
      ('0', "01110110", "0110101100", "0110100011", '0'),
      ('0', "01110111", "1110100011", "0001011100", '1'),
      ('0', "01111000", "1100110011", "0011001100", '1'),
      ('0', "01111001", "1001101100", "1001100011", '0'),
      ('0', "01111010", "0101101100", "0101100011", '0'),
      ('0', "01111011", "1101100011", "0010011100", '1'),
      ('0', "01111100", "0011101100", "0011100011", '0'),
      ('0', "01111101", "1011100011", "0100011100", '1'),
      ('0', "01111110", "0111100011", "1000011100", '1'),
      ('0', "01111111", "1010110011", "0101001100", '1'),
      ('0', "10000000", "1001110010", "0110001101", '0'),
      ('0', "10000001", "0111010010", "1000101101", '0'),
      ('0', "10000010", "1011010010", "0100101101", '0'),
      ('0', "10000011", "1100011101", "1100010010", '1'),
      ('0', "10000100", "1101010010", "0010101101", '0'),
      ('0', "10000101", "1010011101", "1010010010", '1'),
      ('0', "10000110", "0110011101", "0110010010", '1'),
      ('0', "10000111", "1110001101", "0001110010", '1'),
      ('0', "10001000", "1110010010", "0001101101", '0'),
      ('0', "10001001", "1001011101", "1001010010", '1'),
      ('0', "10001010", "0101011101", "0101010010", '1'),
      ('0', "10001011", "1101001101", "1101000010", '1'),
      ('0', "10001100", "0011011101", "0011010010", '1'),
      ('0', "10001101", "1011001101", "1011000010", '1'),
      ('0', "10001110", "0111001101", "0111000010", '1'),
      ('0', "10001111", "0101110010", "1010001101", '0'),
      ('0', "10010000", "0110110010", "1001001101", '0'),
      ('0', "10010001", "1000111101", "1000110010", '1'),
      ('0', "10010010", "0100111101", "0100110010", '1'),
      ('0', "10010011", "1100101101", "1100100010", '1'),
      ('0', "10010100", "0010111101", "0010110010", '1'),
      ('0', "10010101", "1010101101", "1010100010", '1'),
      ('0', "10010110", "0110101101", "0110100010", '1'),
      ('0', "10010111", "1110100010", "0001011101", '0'),
      ('0', "10011000", "1100110010", "0011001101", '0'),
      ('0', "10011001", "1001101101", "1001100010", '1'),
      ('0', "10011010", "0101101101", "0101100010", '1'),
      ('0', "10011011", "1101100010", "0010011101", '0'),
      ('0', "10011100", "0011101101", "0011100010", '1'),
      ('0', "10011101", "1011100010", "0100011101", '0'),
      ('0', "10011110", "0111100010", "1000011101", '0'),
      ('0', "10011111", "1010110010", "0101001101", '0'),
      ('0', "10100000", "1001111010", "0110001010", '1'),
      ('0', "10100001", "0111011010", "1000101010", '1'),
      ('0', "10100010", "1011011010", "0100101010", '1'),
      ('0', "10100011", "1100011010", "1100011010", '0'),
      ('0', "10100100", "1101011010", "0010101010", '1'),
      ('0', "10100101", "1010011010", "1010011010", '0'),
      ('0', "10100110", "0110011010", "0110011010", '0'),
      ('0', "10100111", "1110001010", "0001111010", '0'),
      ('0', "10101000", "1110011010", "0001101010", '1'),
      ('0', "10101001", "1001011010", "1001011010", '0'),
      ('0', "10101010", "0101011010", "0101011010", '0'),
      ('0', "10101011", "1101001010", "1101001010", '0'),
      ('0', "10101100", "0011011010", "0011011010", '0'),
      ('0', "10101101", "1011001010", "1011001010", '0'),
      ('0', "10101110", "0111001010", "0111001010", '0'),
      ('0', "10101111", "0101111010", "1010001010", '1'),
      ('0', "10110000", "0110111010", "1001001010", '1'),
      ('0', "10110001", "1000111010", "1000111010", '0'),
      ('0', "10110010", "0100111010", "0100111010", '0'),
      ('0', "10110011", "1100101010", "1100101010", '0'),
      ('0', "10110100", "0010111010", "0010111010", '0'),
      ('0', "10110101", "1010101010", "1010101010", '0'),
      ('0', "10110110", "0110101010", "0110101010", '0'),
      ('0', "10110111", "1110101010", "0001011010", '1'),
      ('0', "10111000", "1100111010", "0011001010", '1'),
      ('0', "10111001", "1001101010", "1001101010", '0'),
      ('0', "10111010", "0101101010", "0101101010", '0'),
      ('0', "10111011", "1101101010", "0010011010", '1'),
      ('0', "10111100", "0011101010", "0011101010", '0'),
      ('0', "10111101", "1011101010", "0100011010", '1'),
      ('0', "10111110", "0111101010", "1000011010", '1'),
      ('0', "10111111", "1010111010", "0101001010", '1'),
      ('0', "11000000", "1001110110", "0110000110", '1'),
      ('0', "11000001", "0111010110", "1000100110", '1'),
      ('0', "11000010", "1011010110", "0100100110", '1'),
      ('0', "11000011", "1100010110", "1100010110", '0'),
      ('0', "11000100", "1101010110", "0010100110", '1'),
      ('0', "11000101", "1010010110", "1010010110", '0'),
      ('0', "11000110", "0110010110", "0110010110", '0'),
      ('0', "11000111", "1110000110", "0001110110", '0'),
      ('0', "11001000", "1110010110", "0001100110", '1'),
      ('0', "11001001", "1001010110", "1001010110", '0'),
      ('0', "11001010", "0101010110", "0101010110", '0'),
      ('0', "11001011", "1101000110", "1101000110", '0'),
      ('0', "11001100", "0011010110", "0011010110", '0'),
      ('0', "11001101", "1011000110", "1011000110", '0'),
      ('0', "11001110", "0111000110", "0111000110", '0'),
      ('0', "11001111", "0101110110", "1010000110", '1'),
      ('0', "11010000", "0110110110", "1001000110", '1'),
      ('0', "11010001", "1000110110", "1000110110", '0'),
      ('0', "11010010", "0100110110", "0100110110", '0'),
      ('0', "11010011", "1100100110", "1100100110", '0'),
      ('0', "11010100", "0010110110", "0010110110", '0'),
      ('0', "11010101", "1010100110", "1010100110", '0'),
      ('0', "11010110", "0110100110", "0110100110", '0'),
      ('0', "11010111", "1110100110", "0001010110", '1'),
      ('0', "11011000", "1100110110", "0011000110", '1'),
      ('0', "11011001", "1001100110", "1001100110", '0'),
      ('0', "11011010", "0101100110", "0101100110", '0'),
      ('0', "11011011", "1101100110", "0010010110", '1'),
      ('0', "11011100", "0011100110", "0011100110", '0'),
      ('0', "11011101", "1011100110", "0100010110", '1'),
      ('0', "11011110", "0111100110", "1000010110", '1'),
      ('0', "11011111", "1010110110", "0101000110", '1'),
      ('0', "11100000", "1001110001", "0110001110", '0'),
      ('0', "11100001", "0111010001", "1000101110", '0'),
      ('0', "11100010", "1011010001", "0100101110", '0'),
      ('0', "11100011", "1100011110", "1100010001", '1'),
      ('0', "11100100", "1101010001", "0010101110", '0'),
      ('0', "11100101", "1010011110", "1010010001", '1'),
      ('0', "11100110", "0110011110", "0110010001", '1'),
      ('0', "11100111", "1110001110", "0001110001", '1'),
      ('0', "11101000", "1110010001", "0001101110", '0'),
      ('0', "11101001", "1001011110", "1001010001", '1'),
      ('0', "11101010", "0101011110", "0101010001", '1'),
      ('0', "11101011", "1101001110", "1101001000", '1'),
      ('0', "11101100", "0011011110", "0011010001", '1'),
      ('0', "11101101", "1011001110", "1011001000", '1'),
      ('0', "11101110", "0111001110", "0111001000", '1'),
      ('0', "11101111", "0101110001", "1010001110", '0'),
      ('0', "11110000", "0110110001", "1001001110", '0'),
      ('0', "11110001", "1000110111", "1000110001", '1'),
      ('0', "11110010", "0100110111", "0100110001", '1'),
      ('0', "11110011", "1100101110", "1100100001", '1'),
      ('0', "11110100", "0010110111", "0010110001", '1'),
      ('0', "11110101", "1010101110", "1010100001", '1'),
      ('0', "11110110", "0110101110", "0110100001", '1'),
      ('0', "11110111", "1110100001", "0001011110", '0'),
      ('0', "11111000", "1100110001", "0011001110", '0'),
      ('0', "11111001", "1001101110", "1001100001", '1'),
      ('0', "11111010", "0101101110", "0101100001", '1'),
      ('0', "11111011", "1101100001", "0010011110", '0'),
      ('0', "11111100", "0011101110", "0011100001", '1'),
      ('0', "11111101", "1011100001", "0100011110", '0'),
      ('0', "11111110", "0111100001", "1000011110", '0'),
      ('0', "11111111", "1010110001", "0101001110", '0'),
      ('1', "00011100", "0011110100", "1100001011", '0'),
      ('1', "00111100", "0011111001", "1100000110", '1'),
      ('1', "01011100", "0011110101", "1100001010", '1'),
      ('1', "01111100", "0011110011", "1100001100", '1'),
      ('1', "10011100", "0011110010", "1100001101", '0'),
      ('1', "10111100", "0011111010", "1100000101", '1'),
      ('1', "11011100", "0011110110", "1100001001", '1'),
      ('1', "11111100", "0011111000", "1100000111", '0'),
      ('1', "11110111", "1110101000", "0001010111", '0'),
      ('1', "11111011", "1101101000", "0010010111", '0'),
      ('1', "11111101", "1011101000", "0100010111", '0'),
      ('1', "11111110", "0111101000", "1000010111", '0')
    );


end package lookup_8b10b;
